module datamux(
input [15:0] FATECNTR,
input [31:0] FATENDCA,
input [31:0] ERCYBTCNTR,
output reg [7:0] MUXFATBO
);


endmodule 